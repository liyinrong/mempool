`include "common_cells/registers.svh"

module mempool_tile_resp_arbiter #(
    parameter int unsigned NumInp = 16,
    parameter int unsigned AgeMatrixNumEnq = 2,
    parameter int unsigned NumOut = 3,
    parameter type         payload_t   = logic
) (
    input  logic clk_i,
    input  logic rst_ni,

    input  payload_t [NumInp-1:0] data_i,
    input  logic [NumInp-1:0] valid_i,
    output logic [NumInp-1:0] ready_o,

    output payload_t [NumOut-1:0] data_o,
    output logic [NumOut-1:0] valid_o,
    input  logic [NumOut-1:0] ready_i
);

  logic [NumInp-1:0] current_valid_new, current_valid_old;
  logic [NumInp-1:0] current_handshake;

  logic [NumInp-1:0] req_mask_combined_limited_2_new_req; // limit the max new req per cycle to 2

  logic [NumInp-1:0] new_valid_d, new_valid_q, new_valid_d_set, new_valid_d_clr, new_valid_d_en;

  logic [AgeMatrixNumEnq-1:0] enq_fire;
  logic [AgeMatrixNumEnq-1:0] enq_empty;
  logic [AgeMatrixNumEnq-1:0][cf_math_pkg::idx_width(NumInp)-1:0] req_mask_idx;
  logic [AgeMatrixNumEnq-1:0][NumInp-1:0] enq_mask;
  logic [AgeMatrixNumEnq-1:0][NumInp-1:0] req_mask;
  logic [AgeMatrixNumEnq-1:0]             req_mask_vld;
  logic [NumInp-1:0]                      req_mask_combined;

  logic deq_fire;
  logic [NumInp-1:0] deq_mask;

  logic [NumOut-1:0] age_matrix_result_mask_vld;
  logic [NumOut-1:0][NumInp-1:0] age_matrix_result_mask;

  logic [NumOut-1:0] outport_hsk;
  assign outport_hsk = valid_o & ready_i;

  assign current_handshake = valid_i & ready_o;
  assign current_valid_new = valid_i & new_valid_q;
  assign current_valid_old = valid_i & ~new_valid_q;

  // generate the new_valid_q signal, which marks if the valid is new one (which should enqueue age matrix if not hsk) or not
  assign new_valid_d_en   = new_valid_d_set | new_valid_d_clr;
  assign new_valid_d_set  = req_mask_combined_limited_2_new_req & ready_o;
  assign new_valid_d_clr  = req_mask_combined_limited_2_new_req & ~ready_o;
  assign new_valid_d      = (new_valid_q | new_valid_d_set) & ~new_valid_d_clr;

  for (genvar b = 0; b < NumInp; b++) begin
    `FFL(new_valid_q[b], new_valid_d[b], new_valid_d_en[b], '1)
  end

  if(AgeMatrixNumEnq > 2) begin
    $fatal("AgeMatrixNumEnq > 2, this is not supported yet by the age matrix.");
  end

  for (genvar i = 0; i < AgeMatrixNumEnq; i++) begin: gen_enq_fire
    lzc #(
      .WIDTH(NumInp),
      .MODE(i % 2)
    ) i_lzc (
      .in_i(current_valid_new),
      .cnt_o(req_mask_idx[i]),
      .empty_o(enq_empty[i])
    );
    if (i%2 == 0) begin: gen_req_vld_mask_even
      assign req_mask[i] = (1 << req_mask_idx[i]);
    end else begin: gen_req_vld_mask_odd
      logic [NumInp-1:0] req_vld_mask_tmp;
      assign req_vld_mask_tmp = (1 << req_mask_idx[i]);
      for (genvar j = 0; j < NumInp; j++) begin: gen_enq_mask_odd_inner
        assign req_mask[i][j] = req_vld_mask_tmp[NumInp-1 - j];
      end
    end
    assign enq_mask[i] = req_mask[i] & ~current_handshake;

    if (i == 0) begin
      assign req_mask_vld[i]  = ~enq_empty[i];
    end else begin
      assign req_mask_vld[i]  = ~enq_empty[i] & ~(|(req_mask[i] & req_mask[i-1])); // don't choose the same idx as the previous ones
    end
    assign enq_fire[i] = req_mask_vld[i] & |(enq_mask[i]);
  end

  // request shift to let them be mapped to different output ports
  logic [AgeMatrixNumEnq-1:0][NumInp-1:0] req_mask_reordered;
  logic [AgeMatrixNumEnq-1:0]             req_mask_vld_reordered;
  logic [$clog2(AgeMatrixNumEnq)-1:0]     req_mask_reorder_ptr_d, req_mask_reorder_ptr_q;
  assign req_mask_reorder_ptr_d = req_mask_reorder_ptr_q + 1;
  `FFL(req_mask_reorder_ptr_q, req_mask_reorder_ptr_d, 1'b1, '0)

  generate
    if (AgeMatrixNumEnq == 1) begin: gen_req_mask_reorder_1
      assign req_mask_reordered = req_mask;
      assign req_mask_vld_reordered = req_mask_vld;
    end else if (AgeMatrixNumEnq == 2) begin: gen_req_mask_reorder_2
      always_comb begin
        unique case (req_mask_reorder_ptr_q)
          1'b1: begin
            req_mask_reordered[0]  = req_mask[1];
            req_mask_reordered[1]  = req_mask[0];

            req_mask_vld_reordered[0]  = req_mask_vld[1];
            req_mask_vld_reordered[1]  = req_mask_vld[0];
          end
          default: begin
            req_mask_reordered      = req_mask;
            req_mask_vld_reordered  = req_mask_vld;
          end
        endcase
      end
    end else begin: gen_req_mask_reorder_error
      $fatal("AgeMatrixNumEnq > 2, this is not supported yet by the age matrix.");
    end
  endgenerate


  logic [NumOut-1:0][NumInp-1:0] age_matrix_result_mask_reordered;
  logic [NumOut-1:0]             age_matrix_result_mask_vld_reordered;
  logic [$clog2(NumOut)-1:0]     age_matrix_result_mask_reorder_ptr_d, age_matrix_result_mask_reorder_ptr_q;
  assign age_matrix_result_mask_reorder_ptr_d = age_matrix_result_mask_reorder_ptr_q + 1;
  `FFL(age_matrix_result_mask_reorder_ptr_q, age_matrix_result_mask_reorder_ptr_d, 1'b1, '0)

  generate
    if (NumOut == 1) begin: gen_age_matrix_result_mask_reorder_1
      assign age_matrix_result_mask_reordered = age_matrix_result_mask;
      assign age_matrix_result_mask_vld_reordered = age_matrix_result_mask_vld;
    end else if (NumOut == 2) begin: gen_age_matrix_result_mask_reorder_2
      always_comb begin
        unique case (age_matrix_result_mask_reorder_ptr_q)
          1'b1: begin
            age_matrix_result_mask_reordered[0]  = age_matrix_result_mask[1];
            age_matrix_result_mask_reordered[1]  = age_matrix_result_mask[0];

            age_matrix_result_mask_vld_reordered[0]  = age_matrix_result_mask_vld[1];
            age_matrix_result_mask_vld_reordered[1]  = age_matrix_result_mask_vld[0];
          end
          default: begin
            age_matrix_result_mask_reordered      = age_matrix_result_mask;
            age_matrix_result_mask_vld_reordered  = age_matrix_result_mask_vld;
          end
        endcase
      end
    end else if ((NumOut == 3)) begin: gen_age_matrix_result_mask_reorder_3
      always_comb begin
        unique case (age_matrix_result_mask_reorder_ptr_q)
          2'b00: begin
            age_matrix_result_mask_reordered[0]  = age_matrix_result_mask[1];
            age_matrix_result_mask_reordered[1]  = age_matrix_result_mask[2];
            age_matrix_result_mask_reordered[2]  = age_matrix_result_mask[0];

            age_matrix_result_mask_vld_reordered[0]  = age_matrix_result_mask_vld[1];
            age_matrix_result_mask_vld_reordered[1]  = age_matrix_result_mask_vld[2];
            age_matrix_result_mask_vld_reordered[2]  = age_matrix_result_mask_vld[0];
          end
          2'b01: begin
            age_matrix_result_mask_reordered[0]  = age_matrix_result_mask[2];
            age_matrix_result_mask_reordered[1]  = age_matrix_result_mask[0];
            age_matrix_result_mask_reordered[2]  = age_matrix_result_mask[1];

            age_matrix_result_mask_vld_reordered[0]  = age_matrix_result_mask_vld[2];
            age_matrix_result_mask_vld_reordered[1]  = age_matrix_result_mask_vld[0];
            age_matrix_result_mask_vld_reordered[2]  = age_matrix_result_mask_vld[1];
          end
          2'b10: begin
            age_matrix_result_mask_reordered[0]  = age_matrix_result_mask[2];
            age_matrix_result_mask_reordered[1]  = age_matrix_result_mask[1];
            age_matrix_result_mask_reordered[2]  = age_matrix_result_mask[0];

            age_matrix_result_mask_vld_reordered[0]  = age_matrix_result_mask_vld[2];
            age_matrix_result_mask_vld_reordered[1]  = age_matrix_result_mask_vld[1];
            age_matrix_result_mask_vld_reordered[2]  = age_matrix_result_mask_vld[0];
          end
          default: begin
            age_matrix_result_mask_reordered      = age_matrix_result_mask;
            age_matrix_result_mask_vld_reordered  = age_matrix_result_mask_vld;
          end
        endcase
      end
    end else begin: gen_age_matrix_result_mask_reorder_error
      $fatal("NumOut > 3, this is not supported yet by the age matrix.");
    end
  endgenerate

  mux_onehot #(
      .InputWidth(AgeMatrixNumEnq),
      .DataWidth (NumInp)
  ) i_req_mask_combined_mux_onehot (
      .sel_i ('1),
      .data_i(req_mask),
      .data_o(req_mask_combined)
  );

  assign deq_fire = |deq_mask;
  assign deq_mask = current_handshake & ~new_valid_q;

  for (genvar i = 0; i < NumOut; i++) begin: gen_result_mask_vld
    assign age_matrix_result_mask_vld[i] = |age_matrix_result_mask[i];
  end

  age_matrix #(
      .NumEntries (NumInp),
      .NumEnq     (AgeMatrixNumEnq    ),
      .NumSel     (NumOut    )
  ) i_age_matrix (
      .enq_fire_i   (enq_fire           ),
      .enq_mask_i   (enq_mask           ),
      .deq_fire_i   (deq_fire           ),
      .deq_mask_i   (deq_mask           ),
      .sel_mask_i   (current_valid_old  ),
      .result_mask_o(age_matrix_result_mask  ),
      .entry_vld_i  (current_valid_old  ),
      .clk_i        (clk_i              ),
      .rst_ni       (rst_ni             )
  );

  // if agematrix valid output number less than NumOut, choose new request(s) to fit the max output port number
  logic [NumOut+AgeMatrixNumEnq-1:0] combined_mask_valid;
  logic [NumOut+AgeMatrixNumEnq-1:0][NumInp-1:0] combined_mask;

  logic [NumOut-1:0][$clog2(NumOut+AgeMatrixNumEnq)-1:0] sel_inport_idx;
  logic [NumOut-1:0]                                     sel_inport_idx_vld;
  logic [NumOut+AgeMatrixNumEnq-1:0][$clog2(NumOut)-1:0] asn_outport_idx;
  logic [NumOut+AgeMatrixNumEnq-1:0]                     asn_outport_vld;

  assign combined_mask_valid = {req_mask_vld_reordered, age_matrix_result_mask_vld_reordered};
  assign combined_mask       = {req_mask_reordered, age_matrix_result_mask_reordered};

`define ADAPTIVE_REQ_OUTPORT_ALLOC
`ifndef ADAPTIVE_REQ_OUTPORT_ALLOC
  logic [$clog2(NumOut+AgeMatrixNumEnq)-1:0] priority_shift_q, priority_shift_d;
  assign priority_shift_d = priority_shift_q < (NumOut+AgeMatrixNumEnq-1) ? priority_shift_q + 1 : '0;
  `FFL(priority_shift_q, priority_shift_d, 1'b1, '0)
  mempool_tile_resp_select #(
    .InNum  (NumOut+AgeMatrixNumEnq),
    .OutNum (NumOut)
  ) i_mempool_tile_resp_select (
    .req_vector_i         (combined_mask_valid),
    // .priority_i           (priority_shift_q   ),
    .priority_i           ('0 ),
    .sel_inport_idx_o     (sel_inport_idx     ),
    .sel_inport_idx_vld_o (sel_inport_idx_vld ),
    .asn_outport_idx_o    (asn_outport_idx    ),
    .asn_outport_vld_o    (asn_outport_vld    )
  );
`else
  // assign valid requests to ready output ports
  logic [NumOut-1:0][$clog2(NumOut+AgeMatrixNumEnq)-1:0] sel_inport_idx_tmp;
  logic [NumOut-1:0]                                     sel_inport_idx_vld_tmp;
  always_comb begin
    sel_inport_idx_vld_tmp = '0;
    sel_inport_idx_tmp     = '0;
    for (int i = 0; i < (NumOut+AgeMatrixNumEnq); i++) begin
      if (combined_mask_valid[i] == 1'b1) begin
        for (int j = 0; j < NumOut; j++) begin
          if (ready_i[j] == 1'b1) begin
            if (sel_inport_idx_vld_tmp[j] == 1'b0) begin
              sel_inport_idx_tmp[j]     = i;
              sel_inport_idx_vld_tmp[j] = 1'b1;
              break;
            end
          end
        end
      end
    end
  end
  // reorder the output port index to avoid fixed priority
  logic [5-1:0] priority_outport_idx_d, priority_outport_idx_q;
  `FFL(priority_outport_idx_q, priority_outport_idx_d, 1'b1, '0)
  assign priority_outport_idx_d = priority_outport_idx_q < ((1<<5)-1) ? priority_outport_idx_q + 1 : '0;
  if (NumOut == 1) begin: gen_priority_outport_idx_1
    assign sel_inport_idx     = sel_inport_idx_tmp;
    assign sel_inport_idx_vld = sel_inport_idx_vld_tmp;
  end else if (NumOut == 2) begin: gen_priority_outport_idx_2
    always_comb begin
      sel_inport_idx     = '0;
      sel_inport_idx_vld = '0;
      unique case (priority_outport_idx_q[0])
        1'b1: begin
          sel_inport_idx[0]     = sel_inport_idx_tmp[1];
          sel_inport_idx_vld[0] = sel_inport_idx_vld_tmp[1];
          sel_inport_idx[1]     = sel_inport_idx_tmp[0];
          sel_inport_idx_vld[1] = sel_inport_idx_vld_tmp[0];
        end
        default: begin
          sel_inport_idx     = sel_inport_idx_tmp;
          sel_inport_idx_vld = sel_inport_idx_vld_tmp;
        end
      endcase
    end
  end else if (NumOut == 3) begin: gen_priority_outport_idx_3
    localparam int unsigned HASH_BIN = 6; // permutation(NumOut, NumOut)
    logic [5-1:0] hash_out;
    assign hash_out = mempool_pkg::fair_hash(priority_outport_idx_q);
    always_comb begin
      sel_inport_idx     = '0;
      sel_inport_idx_vld = '0;
      unique if ((hash_out >= 0) && (hash_out < HASH_BIN * 1)) begin
        sel_inport_idx[0]     = sel_inport_idx_tmp[0];
        sel_inport_idx_vld[0] = sel_inport_idx_vld_tmp[0];
        sel_inport_idx[1]     = sel_inport_idx_tmp[2];
        sel_inport_idx_vld[1] = sel_inport_idx_vld_tmp[2];
        sel_inport_idx[2]     = sel_inport_idx_tmp[1];
        sel_inport_idx_vld[2] = sel_inport_idx_vld_tmp[1];
      end else if ((hash_out >= HASH_BIN * 1) && (hash_out < HASH_BIN * 2)) begin
        sel_inport_idx[0]     = sel_inport_idx_tmp[1];
        sel_inport_idx_vld[0] = sel_inport_idx_vld_tmp[1];
        sel_inport_idx[1]     = sel_inport_idx_tmp[2];
        sel_inport_idx_vld[1] = sel_inport_idx_vld_tmp[2];
        sel_inport_idx[2]     = sel_inport_idx_tmp[0];
        sel_inport_idx_vld[2] = sel_inport_idx_vld_tmp[0];
      end else if ((hash_out >= HASH_BIN * 2) && (hash_out < HASH_BIN * 3)) begin
        sel_inport_idx[0]     = sel_inport_idx_tmp[2];
        sel_inport_idx_vld[0] = sel_inport_idx_vld_tmp[2];
        sel_inport_idx[1]     = sel_inport_idx_tmp[0];
        sel_inport_idx_vld[1] = sel_inport_idx_vld_tmp[0];
        sel_inport_idx[2]     = sel_inport_idx_tmp[1];
        sel_inport_idx_vld[2] = sel_inport_idx_vld_tmp[1];
      end else if ((hash_out >= HASH_BIN * 3) && (hash_out < HASH_BIN * 4)) begin
        sel_inport_idx[0]     = sel_inport_idx_tmp[2];
        sel_inport_idx_vld[0] = sel_inport_idx_vld_tmp[2];
        sel_inport_idx[1]     = sel_inport_idx_tmp[1];
        sel_inport_idx_vld[1] = sel_inport_idx_vld_tmp[1];
        sel_inport_idx[2]     = sel_inport_idx_tmp[0];
        sel_inport_idx_vld[2] = sel_inport_idx_vld_tmp[0];
      end else if ((hash_out >= HASH_BIN * 4) && (hash_out < HASH_BIN * 5)) begin
        sel_inport_idx[0]     = sel_inport_idx_tmp[1];
        sel_inport_idx_vld[0] = sel_inport_idx_vld_tmp[1];
        sel_inport_idx[1]     = sel_inport_idx_tmp[0];
        sel_inport_idx_vld[1] = sel_inport_idx_vld_tmp[0];
        sel_inport_idx[2]     = sel_inport_idx_tmp[2];
        sel_inport_idx_vld[2] = sel_inport_idx_vld_tmp[2];
      end else begin
        // default case
        sel_inport_idx     = sel_inport_idx_tmp;
        sel_inport_idx_vld = sel_inport_idx_vld_tmp;
      end
      // unique case (priority_outport_idx_q)
      //   2'b00: begin
      //     sel_inport_idx[0]     = sel_inport_idx_tmp[1];
      //     sel_inport_idx_vld[0] = sel_inport_idx_vld_tmp[1];
      //     sel_inport_idx[1]     = sel_inport_idx_tmp[2];
      //     sel_inport_idx_vld[1] = sel_inport_idx_vld_tmp[2];
      //     sel_inport_idx[2]     = sel_inport_idx_tmp[0];
      //     sel_inport_idx_vld[2] = sel_inport_idx_vld_tmp[0];
      //   end
      //   2'b01: begin
      //     sel_inport_idx[0]     = sel_inport_idx_tmp[1];
      //     sel_inport_idx_vld[0] = sel_inport_idx_vld_tmp[1];
      //     sel_inport_idx[1]     = sel_inport_idx_tmp[0];
      //     sel_inport_idx_vld[1] = sel_inport_idx_vld_tmp[0];
      //     sel_inport_idx[2]     = sel_inport_idx_tmp[2];
      //     sel_inport_idx_vld[2] = sel_inport_idx_vld_tmp[2];
      //   end
      //   2'b10: begin
      //     sel_inport_idx[0]     = sel_inport_idx_tmp[1];
      //     sel_inport_idx_vld[0] = sel_inport_idx_vld_tmp[1];
      //     sel_inport_idx[1]     = sel_inport_idx_tmp[2];
      //     sel_inport_idx_vld[1] = sel_inport_idx_vld_tmp[2];
      //     sel_inport_idx[2]     = sel_inport_idx_tmp[0];
      //     sel_inport_idx_vld[2] = sel_inport_idx_vld_tmp[0];
      //   end
      //   default: begin
      //     sel_inport_idx     = sel_inport_idx_tmp;
      //     sel_inport_idx_vld = sel_inport_idx_vld_tmp;
      //   end
      // endcase
    end
  end else begin: gen_priority_outport_idx_error
    $fatal("NumOut > 3, this is not supported yet by the age matrix.");
  end
`endif

  logic [NumOut-1:0][NumInp-1:0] sel_inport_idx_sel_mask;
  logic [NumOut-1:0][$clog2(NumInp)-1:0] sel_inport_idx_sel_mask_bin;
  logic [NumOut-1:0]             sel_inport_idx_sel_mask_vld;
  generate
    for (genvar i = 0; i < NumOut; i++) begin: gen_sel_inport_idx_sel_mask
      assign sel_inport_idx_sel_mask[i]     = combined_mask[sel_inport_idx[i]];
      assign sel_inport_idx_sel_mask_vld[i] = sel_inport_idx_vld[i];

      onehot_to_bin #(
        .ONEHOT_WIDTH   (NumInp)
      ) i_onehot_to_bin (
        .onehot   (sel_inport_idx_sel_mask[i]),
        .bin      (sel_inport_idx_sel_mask_bin[i])
      );
    end
  endgenerate


  assign req_mask_combined_limited_2_new_req = ~(current_valid_new & ~req_mask_combined) & valid_i;


  // data mux
  logic [NumOut-1:0][NumInp-1:0] mux_ready;
  logic [NumInp-1:0][NumOut-1:0] mux_ready_transpose;
  generate
    for (genvar i = 0; i < NumOut; i++) begin: gen_data_mux
      stream_mux #(
        .DATA_T ( payload_t ),
        .N_INP  ( NumInp  )
      ) i_stream_mux (
        .inp_data_i   ( data_i        ),
        .inp_valid_i  ( req_mask_combined_limited_2_new_req & {NumInp{sel_inport_idx_sel_mask_vld[i]}} ),
        .inp_ready_o  ( mux_ready[i]  ),
        .inp_sel_i    ( sel_inport_idx_sel_mask_bin[i] ),
        .oup_data_o   ( data_o[i]     ),
        .oup_valid_o  ( valid_o[i]    ),
        .oup_ready_i  ( ready_i[i]    )
      );
      for (genvar j = 0; j < NumInp; j++) begin: gen_mux_ready_transpose
        assign mux_ready_transpose[j][i] = mux_ready[i][j] & sel_inport_idx_sel_mask_vld[i];
      end
    end 
    for (genvar j = 0; j < NumInp; j++) begin: gen_mux_ready
      assign ready_o[j] = (|mux_ready_transpose[j]) & req_mask_combined_limited_2_new_req[j];
    end
  endgenerate


endmodule
